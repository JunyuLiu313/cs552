/*
   CS/ECE 552 Spring '22
  
   Filename        : memory.v
   Description     : This module contains all components in the Memory stage of the 
                     processor.
*/
`default_nettype none
module memory (/* TODO: Add appropriate inputs/outputs for your memory stage here*/);

   // TODO: Your code here
   
endmodule
`default_nettype wire
