/*
   CS/ECE 552 Spring '22
  
   Filename        : wb.v
   Description     : This is the module for the overall Write Back stage of the processor.
*/
`default_nettype none
module wb (/* TODO: Add appropriate inputs/outputs for your WB stage here*/);

   // TODO: Your code here
   
endmodule
`default_nettype wire
